module video_processor(
	input wire clk_FPGA,   //(50 Mhz)
	input wire clk_en,
	input wire reset,
	input wire [31:0] dataA,
	input wire [31:0] dataB,

	//output wire       done_instruction,
	output wire [2:0] R,
	output wire [2:0] G,
	output wire [2:0] B,
	output wire     out_hsync,
	output wire     out_vsync,
	output reg      out_printtingScreen
);

/*------------------Fios de ligação entre os módulos---------------------*/
wire        new_instruction;
wire 		done;
wire [3:0]  out_opcode;
wire [13:0] out_register;
wire [31:0] out_data;
wire 		done_register;
wire [4:0]  n_reg;
wire [31:0] register_data;
wire 		printtingScreen;
wire [18:0] check_value;
wire [31:0] data_reg;
wire [13:0] memory_address;
wire [13:0] decoded_address;
wire 		active_area;
wire [13:0] address;
wire [8:0]  memory_data;
wire [8:0]  memory_data_out;
wire        done_memory;
wire [8:0]  monitor_color_out;
wire [9:0]  pixel_x;
wire [9:0]  pixel_y;
wire 		clk_100;
wire 		clk_25;
wire        reset_done;
/*------------------------------------------------------------------------*/

/*-----Sinais da unidade de controle para o gerenciamento dos módulos-----*/
wire 	   memory_wr;
//wire [3:0] selectField;
wire 	   register_wr;
wire 	   selectorDemuxRegister;
wire 	   selectorDemuxData;
wire 	   selectorAddress;
wire 	   instruction_finished;
/*------------------------------------------------------------------------*/

reg reg_done;
//reg clk_100;
//reg clk_25;

/*-------Módulo Pll responsável por gerar os sinais de clock necessários para os outros módulos
	c0 - 100 Mhz
	c1 -  25 Mhz
*/

clock_pll clock_pll_inst
(
	.inclk0(clk_FPGA) ,	    // input  inclk0_sig
	.c0(clk_100) ,			// output  c0_sig
	.c1(clk_25) 			// output  c1_sig
);


//background
//32'h3fff1
//32'd12

//sprite
//32'h50
//32'd694310912
decorderInstruction 
decorderInstruction_inst
(
	.clk(clk_100) ,						// input  clk_sig
	.clk_en(clk_en) ,					// input  clk_en_sig
	.dataA(dataA) ,				    // input [31:0] dataA_sig               001010000
	.dataB(dataB) ,				// input [31:0] dataB_sig  101001011000100101100000000000
	.new_instruction(new_instruction) ,	// input  new_instruction_sig
	.out_opcode(out_opcode) ,			// output [1:0]  out_opcode_sig
	.out_register(out_register) ,		// output [13:0] out_register_sig
	.out_data(out_data) 				// output [31:0] out_data_sig
);

controlUnit 
controlUnit_inst
(
	.clk(clk_100) ,							// input  clk_sig
	.reset(!reset) ,							// input  reset_sig
	.opCode(out_opcode) ,					// input [3:0] opCode_sig
	.printtingScreen(printtingScreen) ,		// input  printtingScreen_sig
	.done(instruction_finished) ,			// input  done_sig
	.new_instruction(new_instruction) ,		// output  new_instruction_sig
	.memory_wr(memory_wr) ,					// output  memory_wr_sig
	.selectField() ,						// output [3:0] selectField_sig
	.register_wr(register_wr) ,						// output  register_wr_sig
	.selectorDemuxRegister(selectorDemuxRegister) ,	// output  selectorDemuxRegister_sig
	.selectorDemuxData(selectorDemuxData) ,			// output  selectorDemuxData_sig
	.selectorAddress(selectorAddress), 				// output  selectorAddress_sig
	.reset_done(reset_done)
);


/*--------Demultiplexador para redirecionamento da saída "out_register" do decodificador de instrução--------*/
demultiplexador #(.data_bits(14), .out1_bits_size(14), .out2_bits_size(5), .bits_to_out1(14), .bits_to_out2(5))
demultiplexador_inst_address
(
	.selector(selectorDemuxRegister) ,	// input  selector_sig
	.data(out_register) ,				// input [data_bits-1:0] data_sig
	.out1(decoded_address) ,		    // output [out1_bits_size-1:0] out1_sig (para a memoria)
	.out2(n_reg) 					    // output [out2_bits_size-1:0] out2_sig (para o banco de registradores)
);


/*--------Demultiplexador para redirecionamento da saída "data" do decodificador de instrução--------*/
demultiplexador #(.data_bits(32), .out1_bits_size(9), .out2_bits_size(32), .bits_to_out1(9), .bits_to_out2(32))
demultiplexador_inst_data
(
	.selector(selectorDemuxData) ,		// input  selector_sig
	.data(out_data) ,					// input [data_bits-1:0] data_sig
	.out1(memory_data) ,				// output [out1_bits_size-1:0] out1_sig (para a memoria)
	.out2(register_data) 			    // output [out2_bits_size-1:0] out2_sig (para o banco de registradores)
);


full_register_file full_register_file_inst
(
	.clk(clk_100) ,				// input  clk_sig
	.reset(!reset) ,				// input  reset_sig
	.n_reg(n_reg) ,				// input  n_reg_sig
	.check(check_value) ,		// input [19:0] check_sig
	.written(register_wr) ,		// input  written_sig
	.data(register_data) ,		// input [31:0] data_sig
	.readData(data_reg) ,		// output [31:0] readData_sig
	.success(done_register) 	// output  success_sig
);



full_print_module #(.size_x1(10), .size_y1(10), .size_address1(14), .bits_x_y_1(20), .size_line1(20))
full_print_module_inst
(
	.clk(clk_100) ,								// input  clk_sig
	.clk_pixel(clk_25) ,						// input  clk_pixel_sig
	.reset(!reset) ,								// input  reset_sig
	.data_reg(data_reg) ,						// input [31:0] data_reg_sig
	.active_area(active_area) ,					// input  active_area_sig
	.pixel_x(pixel_x) ,							// input [size_x1-1:0] pixel_x_sig
	.pixel_y(pixel_y) ,							// input [size_y1-1:0] pixel_y_sig
	.memory_address(memory_address) ,	        // output [size_address1-1:0] memory_address_sig
	.printtingScreen(printtingScreen) ,			// output  printtingScreen_sig
	.check_value(check_value) 					// output [bits_x_y_1-1:0] check_value_sig
);

/*-------Multiplexador para selecionar a entrada de endereço para a memória de sprites--------*/
multiplexador #(.data_bits1(14), .data_bits2(14), .out_bits_size(14))
multiplexador_inst
(
	.selector(selectorAddress) ,   	// input  selector_sig
	.data(decoded_address) ,		// input [data_bits1-1:0] data_sig  (vem do decodificador)
	.data2(memory_address) ,		// input [data_bits2-1:0] data2_sig (vem do módulo de impressão)
	.out(address) 					// output [out_bits_size-1:0] out_sig
);

sprite_memory sprite_memory_inst
(
	.address(address) ,					// input [13:0] address_sig
	.clock(clk_100) ,					// input  clock_sig  (100Mhz)
	.reset_done(reset_done),
	.data(memory_data) ,				// input [8:0] data_sig
	.wren(memory_wr) ,					// input  wren_sig
	.out_data(memory_data_out) ,	    // output [8:0] out_data_sig
	.read_memory(done_memory) 	   		// output  read_memory_sig
);


/*------------Módulo para geração do sinais de sincronização do monitor e seus pixeis-----------*/
VGA_sync VGA_sync_inst
(
	.clock(clk_25) ,					// input  clock_sig
	.reset(!reset) ,						// input  reset_sig
	.hsync(out_hsync) ,					// output  hsync_sig
	.vsync(out_vsync) ,					// output  vsync_sig
	.video_enable(active_area) ,	    // output  video_enable_sig
	.pixel_x(pixel_x) ,					// output [9:0] _sig
	.pixel_y(pixel_y) 					// output [8:0] _sig
);

/*
	Bloco combinacional para verificar se um registro no banco de registradores ou uma leitura na memória foi realiza com sucesso.
*/
always @(done_register or done_memory) begin 
	reg_done = done_register | done_memory;
end

/*---------------------Multiplexador que seleciona a saída de cores para o monitor-----------------*/
multiplexador #(.data_bits1(9), .data_bits2(9), .out_bits_size(9))
multiplexador_inst_color
(
	.selector(active_area) ,    // input  selector_sig
	.data(9'b000000000) ,		
	.data2(memory_data_out),    // input [data_bits2-1:0] data2_sig (dados lidos da memória
	.out(monitor_color_out) 	// output [out_bits_size-1:0] out_sig
);


always @(negedge clk_100) begin
	out_printtingScreen  <= printtingScreen;
end

//assign done_instruction = reg_done;
assign instruction_finished = reg_done;
assign R = monitor_color_out[2:0];
assign G = monitor_color_out[5:3];
assign B = monitor_color_out[8:6];

endmodule